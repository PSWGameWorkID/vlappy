module main

fn main() {
	mut i := Game {}
	exit(i.run())
}
